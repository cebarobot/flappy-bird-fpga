`define LCD_5INCH
// `define VGA_640_480
